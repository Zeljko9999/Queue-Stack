`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    15:09:05 06/27/2023 
// Design Name: 
// Module Name:    edge_detector 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module edge_detector(input sig, input clk, output reg edgee);

 reg prethodni_in;

 always@(posedge clk) begin
	prethodni_in <= sig;
	if({prethodni_in, sig} == 2'b01)
		edgee <= 1;
	else
		edgee <= 0;
 end

endmodule